module AvalonBusMaster (

);

endmodule