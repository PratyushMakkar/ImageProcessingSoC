module VGADriver (
  
);
endmodule